`timescale 1ns / 1ps

`include "defines.v"

module mem (
	input wire rst,
	
	// input 
);

endmodule