`timescale 1ns / 1ps

`include "defines.v"

module mem_wb (
	input wire rst,
	input wire clk,
	
	// input 
);

endmodule