`timescale 1ns / 1ps

`include "defines.v"

module wb (
	input wire rst,
	
	// input 
);

endmodule